library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ip_1 is 
    generic (
    );

    port(
    );

end entity;


architecture rtl of ip_1 is

begin

end architecture;


